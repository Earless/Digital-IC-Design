//Verilog HDL for "ICProject", "d_ff_reset" "functional"


module d_ff_reset ( Q, CLK, D, \R~  );

  input \R~ ;
  input CLK;
  input D;
  output Q;
endmodule
